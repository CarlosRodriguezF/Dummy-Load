** Profile: "SCHEMATIC1-Parametrico"  [ C:\Users\Carlos\Documents\DummyLoad\dummy load-pspicefiles\schematic1\parametrico.sim ] 

** Creating circuit file "Parametrico.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "C:\Cadence\SPB_16.5\tools\capture\library\pspice\CSD18502KCS.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
