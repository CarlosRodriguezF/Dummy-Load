** Profile: "SCH-1MOS-Period"  [ C:\Users\Carlos\Documents\DummyLoad\dummy load-pspicefiles\sch-1mos\period.sim ] 

** Creating circuit file "Period.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "C:\Cadence\SPB_16.5\tools\pspice\library\anl_misc.lib" 
.lib "C:\Cadence\SPB_16.5\tools\capture\library\pspice\CSD18502KCS.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 
.STEP PARAM PER LIST 2e-4,5e-5 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCH-1MOS.net" 


.END
